`timescale 1ns/1ps

`define MEM_LIKE_MODULE .clk(clk), .reset(reset),
`define COMB_ONLY_MODULE

`define i(xinstr) data_mem.inner[instr_idx] = xinstr; instr_idx = instr_idx + 1;

module tb_Riscv();
  reg clk, reset;

  wire [31:0] instr_addr;
  wire [31:0] instr;

  wire [31:0] data_addr;
  wire [31:0] mem_read_data;
  wire [31:0] mem_write_data;
  wire should_read_mem;
  wire should_write_mem;

  DataMemory data_mem(`MEM_LIKE_MODULE
    // in
    .instr_addr(instr_addr),
    .data_addr(data_addr),
    .should_write(should_write_mem),
    .write_data(mem_write_data),
    // out
    .instr(instr),
    .read_data(mem_read_data)
  );


  Riscv uut(`MEM_LIKE_MODULE
    // in
    .instr(instr),
    .mem_read_data(mem_read_data),
    // out
    .instr_addr(instr_addr),
    .data_addr(data_addr),
    .should_write_mem(should_write_mem),
    .should_read_mem(should_read_mem),
    .mem_write_data(mem_write_data)
  );

  always #5 clk = ~clk;

  integer instr_idx;
  always @(posedge clk) begin
    // Execute until the instruction memory is out of instructions.
    if (!reset && uut.pc.pc >= instr_idx * 4)
      uut.pc.pc = 0;
  end

  initial begin
    clk = 0;
    reset = 1; #12 reset = 0;
    instr_idx = 0;
    // Initialize the instruction memory with instruction data.

`i(32'h00001137);
`i(32'h00100513);
`i(32'h00100593);
`i(32'h00400613);
`i(32'h00000013);
`i(32'h00000013);
`i(32'h00000013);
`i(32'h00000013);
`i(32'h00000013);
`i(32'h00000097);
`i(32'h000080e7);
`i(32'h0000006f);
`i(32'hfe010113);
`i(32'h00112e23);
`i(32'h00812c23);
`i(32'h00912a23);
`i(32'h01212823);
`i(32'h01312623);
`i(32'h01412423);
`i(32'h00060913);
`i(32'h00058993);
`i(32'h00050413);
`i(32'h00000493);
`i(32'h02600a13);
`i(32'h00040513);
`i(32'h00048593);
`i(32'h00098613);
`i(32'h00090693);
`i(32'h00000097);
`i(32'h000080e7);
`i(32'h00051063);
`i(32'h00148493);
`i(32'h01449063);
`i(32'h00000513);
`i(32'h0000006f);
`i(32'h00100513);
`i(32'h00812a03);
`i(32'h00c12983);
`i(32'h01012903);
`i(32'h01412483);
`i(32'h01812403);
`i(32'h01c12083);
`i(32'h02010113);
`i(32'h00008067);
`i(32'hf3010113);
`i(32'h0c112623);
`i(32'h0c812423);
`i(32'h0c912223);
`i(32'h0d212023);
`i(32'h0b312e23);
`i(32'h0b412c23);
`i(32'h0b512a23);
`i(32'h0b612823);
`i(32'h0b712623);
`i(32'h0b812423);
`i(32'h0b912223);
`i(32'h0ba12023);
`i(32'h09b12e23);
`i(32'h00058793);
`i(32'h02400593);
`i(32'h02b785b3);
`i(32'h00000737);
`i(32'h00070713);
`i(32'h00e585b3);
`i(32'h00c5a107);
`i(32'h0005a007);
`i(32'h0105a187);
`i(32'h0045a087);
`i(32'h5f376737);
`i(32'h9df70b13);
`i(32'h08017253);
`i(32'h0811f1d3);
`i(32'h0145a287);
`i(32'h0085a107);
`i(32'h0185a307);
`i(32'h01c5a587);
`i(32'h0205a607);
`i(32'h0822f553);
`i(32'h080373d3);
`i(32'h0815f353);
`i(32'h082672d3);
`i(32'h106575d3);
`i(32'h1051f653);
`i(32'h08c5f5d3);
`i(32'h10527653);
`i(32'h107576d3);
`i(32'h08d676d3);
`i(32'h1071f653);
`i(32'h10627753);
`i(32'h08e67753);
`i(32'h10b5f653);
`i(32'h10d6f7d3);
`i(32'h00f67653);
`i(32'h000005b7);
`i(32'h00058593);
`i(32'h0005a787);
`i(32'h10e77853);
`i(32'h00c87653);
`i(32'he00605d3);
`i(32'h10f67653);
`i(32'h4015d593);
`i(32'h40bb05b3);
`i(32'hf00587d3);
`i(32'h10f67653);
`i(32'h000005b7);
`i(32'h00058593);
`i(32'h0005a807);
`i(32'h000005b7);
`i(32'h00058593);
`i(32'h0005a887);
`i(32'h10f67653);
`i(32'h01067653);
`i(32'h10f67653);
`i(32'h18c8f7d3);
`i(32'h18f5f653);
`i(32'h18f6f5d3);
`i(32'h00052e87);
`i(32'h00452f07);
`i(32'h00852f87);
`i(32'h18f776d3);
`i(32'h080ef753);
`i(32'h081f77d3);
`i(32'h082ff853);
`i(32'h10c77753);
`i(32'h10b7f7d3);
`i(32'h00f778d3);
`i(32'h00c52707);
`i(32'h01052787);
`i(32'h10d87853);
`i(32'h01187453);
`i(32'h10c77853);
`i(32'h10b7f8d3);
`i(32'h011878d3);
`i(32'h01452807);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052e07);
`i(32'h10d874d3);
`i(32'h0114f8d3);
`i(32'h111474d3);
`i(32'ha09e0553);
`i(32'h00051063);
`i(32'h108774d3);
`i(32'h1087f953);
`i(32'h10887453);
`i(32'h1914f4d3);
`i(32'h19197953);
`i(32'h19147453);
`i(32'h089efed3);
`i(32'h092f7f53);
`i(32'h088fffd3);
`i(32'h080ef4d3);
`i(32'h081f7953);
`i(32'h082fffd3);
`i(32'h10427ed3);
`i(32'h1031ff53);
`i(32'h01eefed3);
`i(32'h10a57f53);
`i(32'h01eeff53);
`i(32'h10727ed3);
`i(32'h1061f453);
`i(32'h008efed3);
`i(32'h10557453);
`i(32'h008efed3);
`i(32'h1073f453);
`i(32'h106379d3);
`i(32'h01347453);
`i(32'h1052f9d3);
`i(32'h013479d3);
`i(32'h10927453);
`i(32'h1121fa53);
`i(32'h01447453);
`i(32'h11f57a53);
`i(32'h008a7453);
`i(32'h1093f4d3);
`i(32'h11237953);
`i(32'h0124f4d3);
`i(32'h11f2ffd3);
`i(32'h009ff953);
`i(32'h113f7fd3);
`i(32'h11def4d3);
`i(32'h089ff4d3);
`i(32'h1089ffd3);
`i(32'h112ef9d3);
`i(32'h093fffd3);
`i(32'h189fffd3);
`i(32'ha1cf95d3);
`i(32'h00000513);
`i(32'h00059063);
`i(32'h112f7e53);
`i(32'h000005b7);
`i(32'h00058593);
`i(32'h0005af07);
`i(32'h108efed3);
`i(32'h09de7e53);
`i(32'h189e7ed3);
`i(32'ha1ee95d3);
`i(32'h00059063);
`i(32'h000005b7);
`i(32'h00058593);
`i(32'h0005ae07);
`i(32'h01dfff53);
`i(32'ha1ee15d3);
`i(32'h00059063);
`i(32'h11f27253);
`i(32'h11f1f1d3);
`i(32'h11f57553);
`i(32'h00407053);
`i(32'h0030f0d3);
`i(32'h00a17153);
`i(32'h11d3f1d3);
`i(32'h11d37253);
`i(32'h11d2f2d3);
`i(32'h0001f353);
`i(32'h001273d3);
`i(32'h0022f553);
`i(32'h00c67053);
`i(32'h00b5f0d3);
`i(32'h00d6f153);
`i(32'h11107053);
`i(32'h1110f0d3);
`i(32'h11117153);
`i(32'h08e07053);
`i(32'h08f0f0d3);
`i(32'h09017153);
`i(32'h200011d3);
`i(32'h20109253);
`i(32'h202112d3);
`i(32'h02612c27);
`i(32'h08612027);
`i(32'h02712a27);
`i(32'h08712227);
`i(32'h02a12827);
`i(32'h08a12427);
`i(32'h10007053);
`i(32'h1010f0d3);
`i(32'h00107053);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052087);
`i(32'h10217153);
`i(32'h00017053);
`i(32'he0000553);
`i(32'h10107053);
`i(32'h40155513);
`i(32'h40ab0533);
`i(32'h000005b7);
`i(32'h00058593);
`i(32'h0005a087);
`i(32'hf0050153);
`i(32'h10207053);
`i(32'h10207053);
`i(32'h00107053);
`i(32'h10207053);
`i(32'h180e7053);
`i(32'h1801f0d3);
`i(32'h08112627);
`i(32'h180270d3);
`i(32'h08112827);
`i(32'h1802f053);
`i(32'h00100513);
`i(32'h08012a27);
`i(32'h00c56063);
`i(32'h00d12023);
`i(32'h00f12223);
`i(32'h00000413);
`i(32'h06012c23);
`i(32'h06012a23);
`i(32'h06012823);
`i(32'h00160493);
`i(32'h08010a13);
`i(32'h07010a93);
`i(32'h02600913);
`i(32'h000a0513);
`i(32'h00040593);
`i(32'h00048613);
`i(32'h000a8693);
`i(32'h00000097);
`i(32'h000080e7);
`i(32'h00051063);
`i(32'h00140413);
`i(32'h01241063);
`i(32'h00000b93);
`i(32'hdeece537);
`i(32'h66d50c13);
`i(32'h00800537);
`i(32'hfff50c93);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052007);
`i(32'h00000d37);
`i(32'h3f000db7);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052087);
`i(32'h02112627);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052087);
`i(32'h02112427);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052087);
`i(32'h02112227);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052087);
`i(32'h02112027);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052087);
`i(32'h00112e27);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052087);
`i(32'h00112c27);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052087);
`i(32'h00112a27);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052087);
`i(32'h00112827);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052087);
`i(32'h00112627);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052087);
`i(32'h00112427);
`i(32'h05810a13);
`i(32'h04810a93);
`i(32'h01000913);
`i(32'h02600993);
`i(32'h02012e27);
`i(32'h04012227);
`i(32'h04012027);
`i(32'h0000006f);
`i(32'h04812007);
`i(32'h04c12087);
`i(32'h05012107);
`i(32'h04412187);
`i(32'h0001f1d3);
`i(32'h04312227);
`i(32'h03c12007);
`i(32'h00107053);
`i(32'h02012e27);
`i(32'h04012007);
`i(32'h00207053);
`i(32'h04012027);
`i(32'h001b8b93);
`i(32'h012b8063);
`i(32'h000d2503);
`i(32'h00000413);
`i(32'h03850533);
`i(32'h00b50513);
`i(32'h019575b3);
`i(32'h01b5e5b3);
`i(32'hf0058053);
`i(32'h03850533);
`i(32'h00b50513);
`i(32'h00ad2023);
`i(32'h01957533);
`i(32'h01b56533);
`i(32'hf00500d3);
`i(32'h10007153);
`i(32'h02c12507);
`i(32'h082571d3);
`i(32'he0018553);
`i(32'h02812587);
`i(32'h10b1f1d3);
`i(32'h40155513);
`i(32'h40ab0533);
`i(32'hf0050253);
`i(32'h1041f1d3);
`i(32'h1041f1d3);
`i(32'h02412607);
`i(32'h083671d3);
`i(32'h1041f1d3);
`i(32'h183571d3);
`i(32'h02012207);
`i(32'h1040f0d3);
`i(32'h1010f253);
`i(32'h1040f2d3);
`i(32'h10527353);
`i(32'h01c12387);
`i(32'h1872f2d3);
`i(32'h0050f0d3);
`i(32'h01812287);
`i(32'h185372d3);
`i(32'h0050f0d3);
`i(32'h104272d3);
`i(32'h10527353);
`i(32'h1052f3d3);
`i(32'h01412687);
`i(32'h10d27253);
`i(32'h00a27253);
`i(32'h01012687);
`i(32'h18d2f2d3);
`i(32'h00527253);
`i(32'h00c12287);
`i(32'h185372d3);
`i(32'h00527253);
`i(32'h00812287);
`i(32'h1853f2d3);
`i(32'h0042f253);
`i(32'h1030f0d3);
`i(32'h103271d3);
`i(32'h03812207);
`i(32'h04412c27);
`i(32'h03412207);
`i(32'h04412e27);
`i(32'h03012207);
`i(32'h06412027);
`i(32'h1010f253);
`i(32'h1031f2d3);
`i(32'h00527253);
`i(32'h00417153);
`i(32'he0010553);
`i(32'h10b17153);
`i(32'h40155513);
`i(32'h40ab0533);
`i(32'hf0050253);
`i(32'h10417153);
`i(32'h10417153);
`i(32'h08267153);
`i(32'h10417153);
`i(32'h18257153);
`i(32'h1820f0d3);
`i(32'h06112227);
`i(32'h1821f0d3);
`i(32'h06112427);
`i(32'h18207053);
`i(32'h06012627);
`i(32'h04012823);
`i(32'h04012623);
`i(32'h04012423);
`i(32'h000a0513);
`i(32'h00040593);
`i(32'h00048613);
`i(32'h000a8693);
`i(32'h00000097);
`i(32'h000080e7);
`i(32'h00051063);
`i(32'h00140413);
`i(32'h01341063);
`i(32'h0000006f);
`i(32'h00000513);
`i(32'h0000006f);
`i(32'h01800513);
`i(32'h02a78533);
`i(32'h000005b7);
`i(32'h00058593);
`i(32'h00a58533);
`i(32'h00c52007);
`i(32'h000005b7);
`i(32'h00058593);
`i(32'h0005a087);
`i(32'h01052107);
`i(32'h01452187);
`i(32'h00107053);
`i(32'h00117153);
`i(32'h0011f0d3);
`i(32'h0006a027);
`i(32'h0026a227);
`i(32'h0016a427);
`i(32'h0000006f);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052007);
`i(32'h04412087);
`i(32'h1000f0d3);
`i(32'h03c12107);
`i(32'h10017153);
`i(32'h07012187);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052207);
`i(32'h07412287);
`i(32'h07812307);
`i(32'h04012387);
`i(32'h1003f053);
`i(32'h1041f1d3);
`i(32'h1042f2d3);
`i(32'h10437253);
`i(32'h0030f0d3);
`i(32'h01800513);
`i(32'h00412583);
`i(32'h02a58533);
`i(32'h000005b7);
`i(32'h00058593);
`i(32'h00b50533);
`i(32'h00052187);
`i(32'h00452307);
`i(32'h00517153);
`i(32'h00407053);
`i(32'h1030f0d3);
`i(32'h10617153);
`i(32'h00852187);
`i(32'h00c52207);
`i(32'h01052287);
`i(32'h01452307);
`i(32'h10307053);
`i(32'h0040f0d3);
`i(32'h00517153);
`i(32'h00607053);
`i(32'h00012503);
`i(32'h00152027);
`i(32'h00252227);
`i(32'h00052427);
`i(32'h00100513);
`i(32'h09c12d83);
`i(32'h0a012d03);
`i(32'h0a412c83);
`i(32'h0a812c03);
`i(32'h0ac12b83);
`i(32'h0b012b03);
`i(32'h0b412a83);
`i(32'h0b812a03);
`i(32'h0bc12983);
`i(32'h0c012903);
`i(32'h0c412483);
`i(32'h0c812403);
`i(32'h0cc12083);
`i(32'h0d010113);
`i(32'h00008067);
`i(32'hfb010113);
`i(32'h04112623);
`i(32'h04812423);
`i(32'h04912223);
`i(32'h05212023);
`i(32'h03312e23);
`i(32'h00000413);
`i(32'hd0157053);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052087);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052107);
`i(32'hd01671d3);
`i(32'h1011f0d3);
`i(32'h18107053);
`i(32'h00207053);
`i(32'hd015f1d3);
`i(32'h1811f0d3);
`i(32'h0020f0d3);
`i(32'h02012027);
`i(32'h02112227);
`i(32'h02012423);
`i(32'h02012623);
`i(32'h02012823);
`i(32'h41200537);
`i(32'h02a12a23);
`i(32'h00012c23);
`i(32'h00012a23);
`i(32'h00012823);
`i(32'h02010913);
`i(32'h01010493);
`i(32'h02600993);
`i(32'h00090513);
`i(32'h00040593);
`i(32'h00000613);
`i(32'h00048693);
`i(32'h00000097);
`i(32'h000080e7);
`i(32'h00051063);
`i(32'h00140413);
`i(32'h01341063);
`i(32'hff000537);
`i(32'h0000006f);
`i(32'h01012007);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052087);
`i(32'h00000537);
`i(32'h00050513);
`i(32'h00052107);
`i(32'h01412187);
`i(32'h28100053);
`i(32'h01812207);
`i(32'h28201053);
`i(32'h281181d3);
`i(32'h282191d3);
`i(32'h00312427);
`i(32'h281200d3);
`i(32'h282090d3);
`i(32'h00112627);
`i(32'he0000553);
`i(32'h00000097);
`i(32'h000080e7);
`i(32'hced91637);
`i(32'h68760413);
`i(32'h40700637);
`i(32'hff760493);
`i(32'h00040613);
`i(32'h00048693);
`i(32'h00000097);
`i(32'h000080e7);
`i(32'h00000097);
`i(32'h000080e7);
`i(32'h00050913);
`i(32'h00812007);
`i(32'he0000553);
`i(32'h00000097);
`i(32'h000080e7);
`i(32'h00040613);
`i(32'h00048693);
`i(32'h00000097);
`i(32'h000080e7);
`i(32'h00000097);
`i(32'h000080e7);
`i(32'h00851993);
`i(32'h00c12007);
`i(32'he0000553);
`i(32'h00000097);
`i(32'h000080e7);
`i(32'h00040613);
`i(32'h00048693);
`i(32'h00000097);
`i(32'h000080e7);
`i(32'h00000097);
`i(32'h000080e7);
`i(32'h01051513);
`i(32'h0129e5b3);
`i(32'h00a5e533);
`i(32'hff0005b7);
`i(32'h00b56533);
`i(32'h03c12983);
`i(32'h04012903);
`i(32'h04412483);
`i(32'h04812403);
`i(32'h04c12083);
`i(32'h05010113);
`i(32'h00008067);
`i(32'hbf000000);
`i(32'h3fc00000);
`i(32'h3f800000);
`i(32'h00000000);
`i(32'h3e4ccccd);
`i(32'h3f000000);
`i(32'h40c90fdb);
`i(32'hc0c00000);
`i(32'h42f00000);
`i(32'hbe800000);
`i(32'h41c00000);
`i(32'hc4340000);
`i(32'h471d8000);
`i(32'h3d800000);
`i(32'h3d23d70a);
`i(32'h3f000000);
`i(32'hbf800000);
`i(32'h3f800000);
`i(32'h00000000);
`i(32'hbeb504f3);
`i(32'hbed2bec2);
`i(32'h3fcb5050);
`i(32'hbf3504f3);
`i(32'hbe257d85);
`i(32'h3fab5050);
`i(32'hbf3504f3);
`i(32'h3e448c60);
`i(32'h3fd8918c);
`i(32'hbeb504f3);
`i(32'hbed2bec2);
`i(32'h3fcb5050);
`i(32'hbf3504f3);
`i(32'h3e448c60);
`i(32'h3fd8918c);
`i(32'hbeb504f3);
`i(32'hbd6dce7c);
`i(32'h3ff8918c);
`i(32'h00000000);
`i(32'hbe257d86);
`i(32'h3fab5050);
`i(32'hbeb504f3);
`i(32'hbed2bec2);
`i(32'h3fcb5050);
`i(32'hbeb504f3);
`i(32'hbd6dce7c);
`i(32'h3ff8918c);
`i(32'h00000000);
`i(32'hbe257d86);
`i(32'h3fab5050);
`i(32'hbeb504f3);
`i(32'hbd6dce7c);
`i(32'h3ff8918c);
`i(32'h00000000);
`i(32'h3e448c5f);
`i(32'h3fd8918c);
`i(32'hbeb504f3);
`i(32'h3db504f2);
`i(32'h3f8b5050);
`i(32'h00000000);
`i(32'hbe257d86);
`i(32'h3fab5050);
`i(32'h00000000);
`i(32'h3e448c5f);
`i(32'h3fd8918c);
`i(32'hbeb504f3);
`i(32'h3db504f2);
`i(32'h3f8b5050);
`i(32'h00000000);
`i(32'h3e448c5f);
`i(32'h3fd8918c);
`i(32'hbeb504f3);
`i(32'h3ee24630);
`i(32'h3fb8918c);
`i(32'hbf3504f3);
`i(32'hbe257d85);
`i(32'h3fab5050);
`i(32'hbeb504f3);
`i(32'h3db504f2);
`i(32'h3f8b5050);
`i(32'hbeb504f3);
`i(32'h3ee24630);
`i(32'h3fb8918c);
`i(32'hbf3504f3);
`i(32'hbe257d85);
`i(32'h3fab5050);
`i(32'hbeb504f3);
`i(32'h3ee24630);
`i(32'h3fb8918c);
`i(32'hbf3504f3);
`i(32'h3e448c60);
`i(32'h3fd8918c);
`i(32'hbf3504f3);
`i(32'h3e448c60);
`i(32'h3fd8918c);
`i(32'hbeb504f3);
`i(32'h3ee24630);
`i(32'h3fb8918c);
`i(32'h00000000);
`i(32'h3e448c5f);
`i(32'h3fd8918c);
`i(32'hbf3504f3);
`i(32'h3e448c60);
`i(32'h3fd8918c);
`i(32'h00000000);
`i(32'h3e448c5f);
`i(32'h3fd8918c);
`i(32'hbeb504f3);
`i(32'hbd6dce7c);
`i(32'h3ff8918c);
`i(32'hbf3504f3);
`i(32'hbe257d85);
`i(32'h3fab5050);
`i(32'hbeb504f3);
`i(32'hbed2bec2);
`i(32'h3fcb5050);
`i(32'h00000000);
`i(32'hbe257d86);
`i(32'h3fab5050);
`i(32'hbf3504f3);
`i(32'hbe257d85);
`i(32'h3fab5050);
`i(32'h00000000);
`i(32'hbe257d86);
`i(32'h3fab5050);
`i(32'hbeb504f3);
`i(32'h3db504f2);
`i(32'h3f8b5050);
`i(32'h3ea7570e);
`i(32'hbf1ffa01);
`i(32'h3f02323a);
`i(32'hbda28f60);
`i(32'hbeba9c88);
`i(32'h3ec14ef0);
`i(32'hbc0dab40);
`i(32'hbd6f5e50);
`i(32'h3f443e88);
`i(32'h3ea7570e);
`i(32'hbf1ffa01);
`i(32'h3f02323a);
`i(32'hbc0dab40);
`i(32'hbd6f5e50);
`i(32'h3f443e88);
`i(32'h3ecb8d8c);
`i(32'hbea34344);
`i(32'h3f65c94a);
`i(32'h3f1c12c1);
`i(32'hbea79fce);
`i(32'h3e647690);
`i(32'h3ea7570e);
`i(32'hbf1ffa01);
`i(32'h3f02323a);
`i(32'h3ecb8d8c);
`i(32'hbea34344);
`i(32'h3f65c94a);
`i(32'h3f1c12c1);
`i(32'hbea79fce);
`i(32'h3e647690);
`i(32'h3ecb8d8c);
`i(32'hbea34344);
`i(32'h3f65c94a);
`i(32'h3f2e2e00);
`i(32'hbcaef100);
`i(32'h3f1cb4b4);
`i(32'h3e505537);
`i(32'hbd892150);
`i(32'h3dbc9710);
`i(32'h3f1c12c1);
`i(32'hbea79fce);
`i(32'h3e647690);
`i(32'h3f2e2e00);
`i(32'hbcaef100);
`i(32'h3f1cb4b4);
`i(32'h3e505537);
`i(32'hbd892150);
`i(32'h3dbc9710);
`i(32'h3f2e2e00);
`i(32'hbcaef100);
`i(32'h3f1cb4b4);
`i(32'h3e8c611a);
`i(32'h3e74d0d4);
`i(32'h3ef653e4);
`i(32'hbda28f60);
`i(32'hbeba9c88);
`i(32'h3ec14ef0);
`i(32'h3e505537);
`i(32'hbd892150);
`i(32'h3dbc9710);
`i(32'h3e8c611a);
`i(32'h3e74d0d4);
`i(32'h3ef653e4);
`i(32'hbda28f60);
`i(32'hbeba9c88);
`i(32'h3ec14ef0);
`i(32'h3e8c611a);
`i(32'h3e74d0d4);
`i(32'h3ef653e4);
`i(32'hbc0dab40);
`i(32'hbd6f5e50);
`i(32'h3f443e88);
`i(32'hbc0dab40);
`i(32'hbd6f5e50);
`i(32'h3f443e88);
`i(32'h3e8c611a);
`i(32'h3e74d0d4);
`i(32'h3ef653e4);
`i(32'h3f2e2e00);
`i(32'hbcaef100);
`i(32'h3f1cb4b4);
`i(32'hbc0dab40);
`i(32'hbd6f5e50);
`i(32'h3f443e88);
`i(32'h3f2e2e00);
`i(32'hbcaef100);
`i(32'h3f1cb4b4);
`i(32'h3ecb8d8c);
`i(32'hbea34344);
`i(32'h3f65c94a);
`i(32'hbda28f60);
`i(32'hbeba9c88);
`i(32'h3ec14ef0);
`i(32'h3ea7570e);
`i(32'hbf1ffa01);
`i(32'h3f02323a);
`i(32'h3f1c12c1);
`i(32'hbea79fce);
`i(32'h3e647690);
`i(32'hbda28f60);
`i(32'hbeba9c88);
`i(32'h3ec14ef0);
`i(32'h3f1c12c1);
`i(32'hbea79fce);
`i(32'h3e647690);
`i(32'h3e505537);
`i(32'hbd892150);
`i(32'h3dbc9710);
`i(32'hbeb504f3);
`i(32'hbf712318);
`i(32'h3f876e74);
`i(32'hbf3504f3);
`i(32'hbf312318);
`i(32'h3f4edce8);
`i(32'hbf3504f3);
`i(32'hbead413c);
`i(32'h3f94afb1);
`i(32'hbeb504f3);
`i(32'hbf712318);
`i(32'h3f876e74);
`i(32'hbf3504f3);
`i(32'hbead413c);
`i(32'h3f94afb1);
`i(32'hbeb504f3);
`i(32'hbf16a09e);
`i(32'h3fb4afb1);
`i(32'h00000000);
`i(32'hbf312318);
`i(32'h3f4edce8);
`i(32'hbeb504f3);
`i(32'hbf712318);
`i(32'h3f876e74);
`i(32'hbeb504f3);
`i(32'hbf16a09e);
`i(32'h3fb4afb1);
`i(32'h00000000);
`i(32'hbf312318);
`i(32'h3f4edce8);
`i(32'hbeb504f3);
`i(32'hbf16a09e);
`i(32'h3fb4afb1);
`i(32'h00000000);
`i(32'hbead413d);
`i(32'h3f94afb1);
`i(32'hbeb504f3);
`i(32'hbee24630);
`i(32'h3f0edce8);
`i(32'h00000000);
`i(32'hbf312318);
`i(32'h3f4edce8);
`i(32'h00000000);
`i(32'hbead413d);
`i(32'h3f94afb1);
`i(32'hbeb504f3);
`i(32'hbee24630);
`i(32'h3f0edce8);
`i(32'h00000000);
`i(32'hbead413d);
`i(32'h3f94afb1);
`i(32'hbeb504f3);
`i(32'hbdb504f4);
`i(32'h3f695f62);
`i(32'hbf3504f3);
`i(32'hbf312318);
`i(32'h3f4edce8);
`i(32'hbeb504f3);
`i(32'hbee24630);
`i(32'h3f0edce8);
`i(32'hbeb504f3);
`i(32'hbdb504f4);
`i(32'h3f695f62);
`i(32'hbf3504f3);
`i(32'hbf312318);
`i(32'h3f4edce8);
`i(32'hbeb504f3);
`i(32'hbdb504f4);
`i(32'h3f695f62);
`i(32'hbf3504f3);
`i(32'hbead413c);
`i(32'h3f94afb1);
`i(32'hbf3504f3);
`i(32'hbead413c);
`i(32'h3f94afb1);
`i(32'hbeb504f3);
`i(32'hbdb504f4);
`i(32'h3f695f62);
`i(32'h00000000);
`i(32'hbead413d);
`i(32'h3f94afb1);
`i(32'hbf3504f3);
`i(32'hbead413c);
`i(32'h3f94afb1);
`i(32'h00000000);
`i(32'hbead413d);
`i(32'h3f94afb1);
`i(32'hbeb504f3);
`i(32'hbf16a09e);
`i(32'h3fb4afb1);
`i(32'hbf3504f3);
`i(32'hbf312318);
`i(32'h3f4edce8);
`i(32'hbeb504f3);
`i(32'hbf712318);
`i(32'h3f876e74);
`i(32'h00000000);
`i(32'hbf312318);
`i(32'h3f4edce8);
`i(32'hbf3504f3);
`i(32'hbf312318);
`i(32'h3f4edce8);
`i(32'h00000000);
`i(32'hbf312318);
`i(32'h3f4edce8);
`i(32'hbeb504f3);
`i(32'hbee24630);
`i(32'h3f0edce8);
`i(32'hc0a9b4a4);
`i(32'h3f07c3b6);
`i(32'h3fc3e1db);
`i(32'h00000000);
`i(32'hc04e0f12);
`i(32'h40a8f876);
`i(32'h40a9b4a4);
`i(32'h3f07c3b6);
`i(32'h3fc3e1db);
`i(32'hc0a9b4a4);
`i(32'h3f07c3b6);
`i(32'h3fc3e1db);
`i(32'h40a9b4a4);
`i(32'h3f07c3b6);
`i(32'h3fc3e1db);
`i(32'h00000000);
`i(32'h4088f876);
`i(32'hc00e0f12);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3f75f5f6);
`i(32'h3f64e4e5);
`i(32'h00000000);
`i(32'h3e888889);
`i(32'h3f64e4e5);
`i(32'h3f6bebec);
`i(32'h3e008081);
`i(32'h3f2dadae);
`i(32'h3f169697);
`i(32'h3e888889);
`i(32'h3f64e4e5);
`i(32'h3f6bebec);
`i(32'h3e008081);
`i(32'h3f2dadae);
`i(32'h3f169697);
`i(32'h3e888889);
`i(32'h3f64e4e5);
`i(32'h3f6bebec);
`i(32'h3e008081);
`i(32'h3f2dadae);
`i(32'h3f169697);
`i(32'h3e888889);
`i(32'h3f64e4e5);
`i(32'h3f6bebec);
`i(32'h3e008081);
`i(32'h3f2dadae);
`i(32'h3f169697);
`i(32'h3e888889);
`i(32'h3f64e4e5);
`i(32'h3f6bebec);
`i(32'h3e008081);
`i(32'h3f2dadae);
`i(32'h3f169697);
`i(32'h3e888889);
`i(32'h3f64e4e5);
`i(32'h3f6bebec);
`i(32'h3e008081);
`i(32'h3f2dadae);
`i(32'h3f169697);
`i(32'h3e888889);
`i(32'h3f64e4e5);
`i(32'h3f6bebec);
`i(32'h3e008081);
`i(32'h3f2dadae);
`i(32'h3f169697);
`i(32'h3e888889);
`i(32'h3f64e4e5);
`i(32'h3f6bebec);
`i(32'h3e008081);
`i(32'h3f2dadae);
`i(32'h3f169697);
`i(32'h3e888889);
`i(32'h3f64e4e5);
`i(32'h3f6bebec);
`i(32'h3e008081);
`i(32'h3f2dadae);
`i(32'h3f169697);
`i(32'h3e888889);
`i(32'h3f64e4e5);
`i(32'h3f6bebec);
`i(32'h3e008081);
`i(32'h3f2dadae);
`i(32'h3f169697);
`i(32'h3e888889);
`i(32'h3f64e4e5);
`i(32'h3f6bebec);
`i(32'h3e008081);
`i(32'h3f2dadae);
`i(32'h3f169697);
`i(32'h3e888889);
`i(32'h3f64e4e5);
`i(32'h3f6bebec);
`i(32'h3e008081);
`i(32'h3f2dadae);
`i(32'h3f169697);
`i(32'h3f66e6e7);
`i(32'h3e48c8c9);
`i(32'h3e8c8c8d);
`i(32'h3f169697);
`i(32'h3e008081);
`i(32'h3e5cdcdd);
`i(32'h3f66e6e7);
`i(32'h3e48c8c9);
`i(32'h3e8c8c8d);
`i(32'h3f169697);
`i(32'h3e008081);
`i(32'h3e5cdcdd);
`i(32'h3f66e6e7);
`i(32'h3e48c8c9);
`i(32'h3e8c8c8d);
`i(32'h3f169697);
`i(32'h3e008081);
`i(32'h3e5cdcdd);
`i(32'h3f66e6e7);
`i(32'h3e48c8c9);
`i(32'h3e8c8c8d);
`i(32'h3f169697);
`i(32'h3e008081);
`i(32'h3e5cdcdd);
`i(32'h3f66e6e7);
`i(32'h3e48c8c9);
`i(32'h3e8c8c8d);
`i(32'h3f169697);
`i(32'h3e008081);
`i(32'h3e5cdcdd);
`i(32'h3f66e6e7);
`i(32'h3e48c8c9);
`i(32'h3e8c8c8d);
`i(32'h3f169697);
`i(32'h3e008081);
`i(32'h3e5cdcdd);
`i(32'h3f66e6e7);
`i(32'h3e48c8c9);
`i(32'h3e8c8c8d);
`i(32'h3f169697);
`i(32'h3e008081);
`i(32'h3e5cdcdd);
`i(32'h3f66e6e7);
`i(32'h3e48c8c9);
`i(32'h3e8c8c8d);
`i(32'h3f169697);
`i(32'h3e008081);
`i(32'h3e5cdcdd);
`i(32'h3f66e6e7);
`i(32'h3e48c8c9);
`i(32'h3e8c8c8d);
`i(32'h3f169697);
`i(32'h3e008081);
`i(32'h3e5cdcdd);
`i(32'h3f66e6e7);
`i(32'h3e48c8c9);
`i(32'h3e8c8c8d);
`i(32'h3f169697);
`i(32'h3e008081);
`i(32'h3e5cdcdd);
`i(32'h3f66e6e7);
`i(32'h3e48c8c9);
`i(32'h3e8c8c8d);
`i(32'h3f169697);
`i(32'h3e008081);
`i(32'h3e5cdcdd);
`i(32'h3f66e6e7);
`i(32'h3e48c8c9);
`i(32'h3e8c8c8d);
`i(32'h3f169697);
`i(32'h3e008081);
`i(32'h3e5cdcdd);
`i(32'h3f800000);
`i(32'h3f800000);
`i(32'h3f800000);
`i(32'h00000000);
`i(32'h00000000);
`i(32'h00000000);

  end

endmodule
